`timescale 1ns/1ns
module row_weight #(parameter M=8,
                    parameter S=8,
                    parameter n=32,
                    parameter cl=8,
                    parameter addrwidth=2)(
        input [addrwidth:0] addr,
        output [M*(n+cl)-1 : 0] W
);

    reg [M*(n+cl)-1 : 0] weight[S:0] ;
    initial begin
        weight[0]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[1]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[2]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[3]={24'h106600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[4]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[5]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[6]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[7]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[8]='b0;
    #63;
        weight[0]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[1]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[2]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[3]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[4]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[5]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[6]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[7]={24'h006600,24'h006600,24'h806689,24'h006600,24'h806689,24'h806689,24'h006600,24'h006600};
        weight[8]='b0;
        /*weight[0]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[1]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[2]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[3]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[4]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[5]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[6]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};
        weight[7]={16'h0066,16'h0066,16'h8066,16'h0066,16'h8066,16'h8066,16'h0200,16'h0200};*/
    end

assign W = weight[addr];

endmodule