library verilog;
use verilog.vl_types.all;
entity tb_row_weight is
end tb_row_weight;
