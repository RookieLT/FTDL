library verilog;
use verilog.vl_types.all;
entity tb_crc is
end tb_crc;
