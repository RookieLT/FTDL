library verilog;
use verilog.vl_types.all;
entity tb_adder_tree is
end tb_adder_tree;
