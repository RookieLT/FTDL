library verilog;
use verilog.vl_types.all;
entity tb_tmr_adder_tree is
end tb_tmr_adder_tree;
