library verilog;
use verilog.vl_types.all;
entity tb_rmac is
end tb_rmac;
