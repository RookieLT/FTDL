library verilog;
use verilog.vl_types.all;
entity tb_tmr_multiplier is
end tb_tmr_multiplier;
