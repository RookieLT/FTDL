library verilog;
use verilog.vl_types.all;
entity tb_ctrl is
end tb_ctrl;
