library verilog;
use verilog.vl_types.all;
entity tb_s2neuron is
end tb_s2neuron;
