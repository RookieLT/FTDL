`timescale 1ns/1ns
module column_weight #(parameter N=8,
                    parameter S=8,
                    parameter n=32,
                    parameter cl=8,
                    parameter addrwidth=2)(
        input [addrwidth:0] addr,
        //output [N*n-1 : 0] W
        output [N*(n+cl)-1 : 0] W
);


    reg [N*(n+cl)-1 : 0] weight[S:0] ;
    //reg [N*n-1 : 0] weight[S-1:0] ;
    initial begin
       
        weight[0]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[1]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[2]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[3]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[4]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[5]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[6]={24'h940095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[7]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[8]='b0;
        #111;
         weight[0]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[1]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[2]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[3]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[4]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[5]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[6]={24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095,24'h840095};
        weight[7]={24'h04001c,24'h04001c,24'h04001c,24'h04001c,24'h04ff1c,24'h04001c,24'h04001c,24'h04001c};
        weight[8]='b0;
        /*
        weight[0]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[1]={16'h0400,16'h0400,16'h0400,16'h0400,16'h04ff,16'h0400,16'h0400,16'h0400};
        weight[2]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[3]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        weight[4]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[5]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        weight[6]={16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400,16'h8400};
        weight[7]={16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400,16'h0400};
        */
    end

assign W = weight[addr];

endmodule